//***************************************************
//*   Регистры видеоконтроллера
//*************************************************
module vregs 
 #(parameter SPEED=19200) // начальная скорость интерфейса по умолчанию
(
// шина wishbone
   input                  wb_clk_i,   // тактовая частота шины
   input                  wb_rst_i,   // сброс
   input    [15:0]        wb_adr_i,   // адрес 
   input    [15:0]        wb_dat_i,   // входные данные
   output reg [15:0]      wb_dat_o,   // выходные данные
   input                  wb_cyc_i,   // начало цикла шины
   input                  wb_we_i,    // разрешение записи (0 - чтение)
   input                  wb_stb_i,   // строб цикла шины
   input    [1:0]         wb_sel_i,   // выбор конкретных байтов для записи - старший, младший или оба
   output reg             wb_ack_o,   // подтверждение выбора устройства
   
   input  [2:0]          initspeed,   // начальная скорость последовательного порта - запишется в регистр конфигурации
// регистры 
   output reg [12:0]     cursor,      // регистр адреса курсора, base+0
   output reg [15:0]     vtcsr        // управляющий регистр,    base+2
);
//-----------------------------------------------------------------------------------------------------
//  base+0  регистр адреса курсора, содержит абсолютный адрес байта с курсором в области видеопамяти
//-----------------------------------------------------------------------------------------------------
//  base+2   Регистр управления терминалом VTCSR:
//  
//   D0: 0 - локальная петля, 1 - связь с ЭВМ
//   D1: 
//   D2: 0 - курсор невидим, 1 - отображается
//   D3: форма курсора: 0 - подчеркивание, 1 - блок
//   D4: 1 - звуковой сигнал
//   D5: импульсы управления мерцанием знаков (0 - знак погашен, 1 - отображается)
//
//   D8..D10: скорость интерфейса:
//            000 - 1200
//            001 - 2400
//            010 - 4800
//            011 - 9600
//            100 - 19200
//            101 - 38400
//            110 - 57600
//            111 - 115200

wire bus_strobe;          // строб шинной транзакции
wire re;                  // строб чтения
wire we;                  // строб записи четных байтов
wire wo;                  // строб записи нечетных байтов

//****************************************   
// Сигналы запроса доступа от шины
//****************************************   
// строб цикла шины
assign bus_strobe = wb_cyc_i & wb_stb_i;         
// чтение
assign re = bus_strobe & ~wb_we_i; 
// запись четных байтов
assign we = bus_strobe & wb_we_i & wb_sel_i[0];
// запись нечетных байтов
assign wo = bus_strobe & wb_we_i & wb_sel_i[1];
// формирователь ответа на цикл шины   
wire reply=wb_cyc_i & wb_stb_i & ~wb_ack_o;
// Сигнал ответа 
always @(posedge wb_clk_i or posedge wb_rst_i)
   if (wb_rst_i == 1'b1) wb_ack_o <= 1'b0;
   else wb_ack_o <= reply;

//****************************************   
//*  Обработка транзакций общей шины
//****************************************   
always @(posedge wb_clk_i or posedge wb_rst_i)
   // сброс
   if (wb_rst_i == 1'b1) begin
       cursor <= {13{1'b0}} ;   // курсор в позиции 0
       vtcsr <= {5'b0000, initspeed,8'b00001};  // сразу включается режим online, устанавливаем скорость по умолчанию
   end   
         
   else begin
       if (re == 1'b1) begin
         // чтение регистров
           if (wb_adr_i[1])  wb_dat_o <= vtcsr;  // регистр управления
          // else wb_dat_o <= {3'b000, cursor} ; // регистр курсора - чтение не требуется
       end 
       else begin
       // запись регистров
          if (wo == 1'b1)   
          // запись нечетных байтов
                if (wb_adr_i[1] == 0) cursor[12:8] <= wb_dat_i[12:8] ;  // регистр курсора
                else vtcsr[15:8] <= wb_dat_i[15:8];  // регистр управления 
               
          if (we == 1'b1)  
             // запись четных байтов 
               if (wb_adr_i[1] == 0) cursor[7:0] <= wb_dat_i[7:0] ; // регистр курсора        
               else vtcsr[7:0] <= wb_dat_i[7:0];  // регистр управления    
             end 
   end 
endmodule
